---------------------------------------------------------------------------------------------------
--
-- Title       : ordenar_extSigno
-- Design      : tipo_b
-- Author      : mario
-- Company     : UTM
--
---------------------------------------------------------------------------------------------------
--
-- File        : C:\My_Designs\procesadorB\tipo_b\compile\ordenar_extSigno.vhd
-- Generated   : Tue Jan 14 22:04:35 2025
-- From        : C:\My_Designs\procesadorB\tipo_b\src\ordenar_extSigno.bde
-- By          : Bde2Vhdl ver. 2.6
--
---------------------------------------------------------------------------------------------------
--
-- Description : 
--
---------------------------------------------------------------------------------------------------
-- Design unit header --
library IEEE;
use IEEE.std_logic_1164.all;


entity ordenar_extSigno is
  port(
       fun7 : in STD_LOGIC_VECTOR(6 downto 0);
       rd : in STD_LOGIC_VECTOR(4 downto 0);
       salida_ordenada : out STD_LOGIC_VECTOR(11 downto 0)
  );
end ordenar_extSigno;

architecture ordenar_extSigno of ordenar_extSigno is

begin

end ordenar_extSigno;

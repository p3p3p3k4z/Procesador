library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL; 

entity memoria_del_programa is
    Port (
        a   : in STD_LOGIC_VECTOR(11 downto 0); -- Entrada del contador de programa (5 bits)
        do  : out STD_LOGIC_VECTOR(31 downto 0) -- Salida de bits de instrucci�n
    );
end memoria_del_programa;

architecture Behavioral of memoria_del_programa is

    type mem_array is array (0 to 60) of STD_LOGIC_VECTOR(31 downto 0);
    
    signal memInstr : mem_array := (
        0 => "00000101100100000000010100010011",-- add x19,x21,x20--"00000000001000011000010100110011", -- ADD
        1 => "00000000001000011000010100010011", -- ADDI  
        2 => "00000000010010011010101100000011", -- lw 
        3 => "11111111111111111111111111111111", 
        4 => "00000011011100000000010110010011", --"11111111111010011000101010010011",-- addi x21,x19,-2 --"01000000001000011000010100110011", -- SUB 
        5 => "11111111111000011000010100010011", -- ADD NEG 
        6 => "00000000011100100010010000100011", -- sw
        7 => "00001111000011110000111100001111", 
        8 => "00000000101000100010000000100011",-- lw x21, 4(x20 --"00000000001000011111010100110011", -- AND 
        9 => "00000000001000011111010100010011", -- ANDI
        10 => "00000000000000000000000000000000", -- nada apartir
        11 => "00001111000011110000111100001111", 
        12 => "00000000101101000010000000100011",-- sw x19, 8(x20) --"00000000001000011110010100110011", -- OR 
        13 => "00000000001000011110010100010011", -- ORI
        14 => "00000000000000000000000000000000", -- lbu
        15 => "00000000000011110000000000001111",
        16 => "00000100101100000000000001100011",--"00000000100000000010101010000011",-- lw x21, 8(x0) --"00000000001000011100010100110011", -- XOR
        17 => "00000000001000011100010100010011", -- XORI
        18 => "00000000000000000000000000000000", -- lhu
        19 => "11111111111111111010101010101010",
        20 => "00000000000001010000011110010011", -- STL
        21 => "00000000001000011010010100010011", -- STLI
        22 => "00000000000000000000000000000000", -- sb
        23 => "11111111111100001111000011110000",
        24 => "00000000101101111100110001100011",-- "00000000001000011011010100110011", -- STLU
        25 => "00000000001000011011010100010011", -- STLUI
        26 => "00000000000000000000000000000000", -- sh
        27 => "11110000000000000000111111111111",
        28 => "01000000101101111000011110110011",-- SLL
        29 => "00000000001000011001010100010011",-- SLLI
        30 => "00000000000000000000000000000000",-- sw
        31 => "00000000000000000000000000000000",
		32 => "11111110111100000001100011100011", -- SRL
		33 => "00000000001000011101010100010011", -- SRLI
		34 => "00000000000000000000000000000000", -- nada
		35 => "11111111111111111111111111111111",
		36 => "00000000000001011000010100010011", -- SRLA 
		37 => "01000000001000011101010100010011", -- SRLAI
		38 => "00000000000000000000000000000000",  -- nada
		39 => "00000000000000000000000000000000",
		40 => "00000000000001111000010110010011",
		41 => "00000000000000000000000000000000",
		42 => "00000000000000000000000000000000",
		43 => "00000000000000000000000000000000",
		44 => "11111010000000000000110011100011",
		45 => "00000000000000000000000000000000",
		46 => "00000000000000000000000000000000",
		47 => "00000000000000000000000000000000",
		48 => "00000000101000000010000000100011",
		49 => "00000000000000000000000000000000",
		50 => "00000000000000000000000000000000",
		51 => "00000000000000000000000000000000",
		52 => "00000000000001010000111100010011",
		53 => "00000000000000000000000000000000",
		54 => "00000000000000000000000000000000",
		55 => "00000000000000000000000000000000",
		56 => "00000000000000000000000001100011",
		57 => "00000000000000000000000000000000",
		58 => "00000000000000000000000000000000",
		59 => "00000000000000000000000000000000",
		60 => "00000000000000000000000000000000"
    );
begin

    do <= memInstr(conv_integer(a)); 
    
end Behavioral;
